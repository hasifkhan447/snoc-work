name=NMOS_PMOS_SWEEP only_toplevel=true spice_ignore=false value="
.options savecurrents

.control
save all

setplot const
let nmos_index = 0
let nmos_w = 10
let nmos_final = 20 
let nmos_step = 1

let nmos_length = ceil((nmos_final - nmos_w)/nmos_step)

let pmos_initial = nmos_w
let pmos_w = pmos_initial
let pmos_final = 40
let pmos_step = 1

let switching_points = vector(nmos_length)
let asymmetricity = vector(nmos_length)
let Rdon_pmos = vector(nmos_length)
let Rdon_nmos = vector(nmos_length)
let rise_times = vector(nmos_length)
let fall_times = vector(nmos_length)
let propagation_delay = vector(nmos_length)
let ratio = vector(nmos_length)
let nmos_width = vector(nmos_length)

set tranplots = ' '
set swplots = ' '

while nmos_w < nmos_final 

  alter m.xm1.msky130_fd_pr__nfet_01v8 W = nmos_w
  alter m.xm3.msky130_fd_pr__nfet_01v8 W = e *nmos_w
  alter m.xm5.msky130_fd_pr__nfet_01v8 W = e * e * nmos_w


  let minimum_delay = 100
  let minimum_width_pmos = 100

  let pmos_w = pmos_initial

**** Find least asymmetric pmos_w **** 
  while pmos_w < pmos_final

    alter m.xm2.msky130_fd_pr__pfet_01v8 W = pmos_w
    alter m.xm4.msky130_fd_pr__pfet_01v8 W = e * pmos_w
    alter m.xm4.msky130_fd_pr__pfet_01v8 W = e * e * pmos_w

* Run transient analysis using a symmetric pulse of period 25n
    tran 10p 40n 

    meas tran rise_time TRIG v(out) VAL=0.1 RISE=LAST TARG v(out) VAL=1.62 RISE=LAST
    meas tran fall_time TRIG v(out) VAL=1.62 FALL=1 TARG v(out) VAL=0.1 FALL=1
* Create array of diffs
    let prop_delay = ( $&rise_time + $&fall_time )/2

    if prop_delay < minimum_delay
      let minimum_delay = prop_delay       
      let minimum_width_pmos = pmos_w
    end
    print prop_delay prop_delay minimum_width_pmos pmos_w
    print nmos_w pmos_w
    let pmos_w = pmos_w + pmos_step
  end

  alter m.xm2.msky130_fd_pr__pfet_01v8 W = minimum_width_pmos
  alter m.xm4.msky130_fd_pr__pfet_01v8 W = e *minimum_width_pmos
  alter m.xm6.msky130_fd_pr__pfet_01v8 W = e * e * minimum_width_pmos


**** Run trainsient again to get rise fall time ****
  tran 10p 40n 
*** Second rise because transient artifacts are technically rises and falls
  meas tran tau_rise TRIG v(out) VAL=0 RISE=LAST TARG v(out) VAL=1.376 RISE=LAST
  meas tran tau_fall TRIG v(out) VAL=1.8 FALL=1 TARG v(out) VAL=0.6624 FALL=1


  let Rdon_nmos[nmos_index] = tau_fall/200f
  let Rdon_pmos[nmos_index] = tau_rise/200f
  let propagation_delay[nmos_index] = minimum_delay

  set tranplots = ( $tranplots {$curplot}.v(out) )

**** Find switching point for aforementioned pmos_w ****

  dc vin 0 1.8 1m 

  meas dc switching_point WHEN v(out)=0.9 CROSS=1

  let switching_points[nmos_index] = $&switching_point
  let ratio[nmos_index] = minimum_width_pmos/nmos_w
  let nmos_width[nmos_index] = nmos_w 
  let propagation_delay[nmos_index] = minimum_delay
  print nmos_index minimum_width_pmos 

  set swplots = ( $swplots {$curplot}.v(out) )


  let nmos_w = nmos_w + nmos_step
  let nmos_index = nmos_index + 1
end

set swplots = ( $swplots {$curplot}.v(in) )

plot switching_points vs ratio xlabel 'W_p/W_n' ylabel 'Switching point' pointplot 
plot Rdon_pmos Rdon_nmos vs ratio xlabel 'W_p/W_n' ylabel 'R_don' pointplot 
plot propagation_delay vs ratio  xlabel 'W_p/W_n' ylabel 'Propagation delay' pointplot 
plot ratio vs nmos_w xlabel 'W_n' ylabel 'W_p/W_n' pointplot 

set nolegend

*plot $swplots xlimit 800m 1 title 'Switching point envelope' 
*plot $tranplots xlimit 1n 3n title 'Transient fall envelope'
*plot $tranplots xlimit 26n 28n title 'Transient rise envelope'


.endc
"










