name=STIMULUS1 only_toplevel=true spice_ignore=false value="
.options savecurrents

.control
save all

let step=1
let final_w_pmos=80
let current_w_pmos=10

let total_iterations = ceil((final_w_pmos - current_w_pmos)/step)
let index= 0

let switching_points = vector(total_iterations)
let asymmetricity = vector(total_iterations)
let width = vector(total_iterations)


while current_w_pmos < final_w_pmos

	alter m.xm2.msky130_fd_pr__pfet_01v8 W=current_w_pmos

******* Asymmetricity analysis ********
	tran 10p 50n ; Run transient analysis using a symmetric pulse of period 25n

	meas tran rise_time TRIG v(out) VAL=0.1 RISE=1 TARG v(out) VAL=1.62 RISE=1 
	meas tran fall_time TRIG v(out) VAL=1.62 FALL=1 TARG v(out) VAL=0.1 FALL=1
	
	let asymmetricity[index] = abs( $&rise_time - $&fall_time ) ; Create array of diffs



******* Switching point analysis ********
	dc vin 0 1.8 1m ; Run dc analysis, check for operating point

	meas dc switching_point WHEN v(out)=v(in) CROSS=LAST
	set plotstr = ( $plotstr {$curplot}.v(out) )  
	set global_switching_point = $&switching_point

	let switching_points[index] = $&switching_point
	let width[index] = current_w_pmos


	let current_w_pmos=current_w_pmos + step
	let index=index + 1

	end

set plotstr = ( $plotstr {$curplot}.v(in) )

set nolegend

******* Plot results ********
plot switching_points vs width title 'switching points vs time' xlabel 'width' ylabel 'Switching point (V)'
plot asymmetricity vs width title 'asymmetricity vs time' xlabel 'width' ylabel 'Difference in rise/fall'

plot $plotstr

******* Find switching point at most symmetric w ********
let lowest_asym = 100
let best_w_index = 0 ; Find most symmetric w
let index = 0
let tolerance = 1p ; We let the asymmetricity be plus/minus 1p of 0 

repeat $&total_iterations 

  let asym = abs(asymmetricity[index] - 1p)
  let current_w_pmos = width[index]

  if asym < lowest_asym ; If we have something smaller, set it as the best goal and repeat
    let best_w_index = index
    let lowest_asym = asym

  end
  
  let index = index + 1
end

* Now that we have the best width, we now need to move towards getting the switching point

let chosen_switching_point = switching_points[best_w_index]
print chosen_switching_point

.endc
"




