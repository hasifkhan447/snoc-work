name=FIXED_NMOS only_toplevel=true spice_ignore=false value="
.options savecurrents

.control
save all

setplot const
let net_switching_points = vector(5)
let nmos_index = 0

set nmos_vals = ( 10 20 30 )
set pmos_vals = ( 10 20 30 )
set length_nmos_vals = 3
set length_pmos_vals = 3

foreach nmos_w $nmos_vals

  alter @m.xm1.msky130_fd_pr__nfet_01v8[w]=nmos_w

  setplot const
  let switching_points = vector($length_nmos_vals)
  let asymmetricity = vector($length_nmos_vals)
  let width = vector($length_nmos_vals)

  let minimum = 100
  set minimum_index = 0

  let index = 0

**** Find least asymmetric pmos_w **** 
  foreach pmos_w $pmos_vals

    alter @m.xm2.msky130_fd_pr__pfet_01v8[w] = pmos_w

  ******* Asymmetricity analysis ********
    tran 10p 50n ; Run transient analysis using a symmetric pulse of period 25n

    meas tran rise_time TRIG v(out) VAL=0.1 RISE=1 TARG v(out) VAL=1.62 RISE=1 
    meas tran fall_time TRIG v(out) VAL=1.62 FALL=1 TARG v(out) VAL=0.1 FALL=1
    
    let diff = abs( $&rise_time - $&fall_time ) ; Create array of diffs

    if diff < minimum
      let minimum = diff       
      let minimum_index = index
    end
    let index = index + 1
  end

  alter @m.xm2.msky130_fd_pr__pfet_01v8[W] = $pmos_vals[minimum_index]

**** Find switching point for aforementioned pmos_w ****

  dc vin 0 1.8 1m ; Run dc analysis, check for operating point

  meas dc switching_point WHEN v(out)=v(in) CROSS=LAST

  let switching_points[nmos_index] = $&switching_point
  let width[nmos_index] = $nmos_w
  let nmos_index = nmos_index + 1
 

end

plot switching_points vs width

.endc
"
