name=VARY_NMOS only_toplevel=true spice_ignore=false value="
*.options savecurrents

.control

setplot new 
set nmos = $curplot
set curplotname = nmos

let step_nmos=1
let index_nmos=0
let final_w_nmos=11
let current_w_nmos=10



let total_iterations_nmos = ceil((final_w_nmos - current_w_nmos)/step_nmos)

setplot new 
set final = $curplot
set curplotname = final

let width_nmos = vector({$nmos}.total_iterations_nmos)
let width_pmos = vector({$nmos}.total_iterations_nmos)
let switching_points = vector({$nmos}.total_iterations_nmos)
let asym = vector({$nmos}.total_iterations_nmos)

setplot new 
set pmos = $curplot
set curplotname = pmos

let current_w_pmos=10

let lowest_asym = 100
let best_w_pmos = 0 


let step_pmos=1
let index_pmos= 0
let final_w_pmos=30



set curplot = $nmos
***** Start varying nmos widths ****
while current_w_nmos < final_w_nmos
  alter @m.xm1.msky130_fd_pr__nfet_01v8[w]=current_w_nmos

* new plot for pmos
  set curplot = $pmos


**** Start varying pmos widths ******
  while current_w_pmos < final_w_pmos

* Set pmos
    alter @m.xm2.msky130_fd_pr__pfet_01v8[w]=current_w_pmos
******* Asymmetricity simulation with pulse of 50n with 1/2 duty cycle ********
    tran 10p 50n 

    meas tran rise_time TRIG v(out) VAL=0.1 RISE=1 TARG v(out) VAL=1.62 RISE=1 
    meas tran fall_time TRIG v(out) VAL=1.62 FALL=1 TARG v(out) VAL=0.1 FALL=1
    let difference = abs( $&rise_time - $&fall_time ) 

    let current_minimum = {$pmos}.lowest_asym
    let current_width = {$pmos}.current_w_pmos

    set aux = $curplot

    if difference < current_minimum
      setplot $pmos
      let lowest_asym = {$aux}.difference 
      let best_w_pmos = current_width
    end
  end 


******* Get switching point of best width ********
  alter m.xm2.msky130_fd_pr__pfet_01v8 W= {$pmos}.best_w_pmos

  dc vin 0 1.8 1m 

  meas dc switching_point WHEN v(out)=v(in) CROSS=LAST

  set aux = $curplot
  setplot $final

  let switching_points[{$pmos}.index_pmos] = {$aux}.switching_point
  let width_pmos[{$pmos}.index_pmos] = {$pmos}.current_w_pmos
  let asym[{$pmos}.index_pmos] = {$pmos}.lowest_asym 

  setplot $nmos
  let index_nmos = index_nmos + 1
  let current_w_nmos = current_w_nmos + step_nmos

end

**** Stop varying nmos widths **** 

set nolegend

******* Plot results ********
plot {$final}.switching_points vs {$final}.width_nmos
plot {$final}.asym vs {$final}.width_nmos
.endc
"

name=FIXED_NMOS only_toplevel=true spice_ignore=false value="
.options savecurrents

.control
save all

foreach nmos_w 10 20 
  alter @m.xm1.msky130_fd_pr__nfet_01v8[w]=$nmos_w

  let step=1
  let final_w_pmos=80
  let current_w_pmos=10

  let total_iterations = ceil((final_w_pmos - current_w_pmos)/step)
  let index= 0

  let switching_points = vector(total_iterations)
  let asymmetricity = vector(total_iterations)
  let width = vector(total_iterations)


  while current_w_pmos < final_w_pmos

    alter m.xm2.msky130_fd_pr__pfet_01v8 W=current_w_pmos

  ******* Asymmetricity analysis ********
    tran 10p 50n ; Run transient analysis using a symmetric pulse of period 25n

    meas tran rise_time TRIG v(out) VAL=0.1 RISE=1 TARG v(out) VAL=1.62 RISE=1 
    meas tran fall_time TRIG v(out) VAL=1.62 FALL=1 TARG v(out) VAL=0.1 FALL=1
    
    let asymmetricity[index] = abs( $&rise_time - $&fall_time ) ; Create array of diffs



  ******* Switching point analysis ********
    dc vin 0 1.8 1m ; Run dc analysis, check for operating point

    meas dc switching_point WHEN v(out)=v(in) CROSS=LAST
    set plotstr = ( $plotstr \{$curplot\}.v(out) )  
    set global_switching_point = $&switching_point

    let switching_points[index] = $&switching_point
    let width[index] = current_w_pmos


    let current_w_pmos=current_w_pmos + step
    let index=index + 1

  end

  set plotstr = ( $plotstr \{$curplot\}.v(in) )

  set nolegend

  ******* Plot results ********
  plot switching_points vs width title 'switching points vs time' xlabel 'width' ylabel 'Switching point (V)'
  plot asymmetricity vs width title 'asymmetricity vs time' xlabel 'width' ylabel 'Difference in rise/fall'

  plot $plotstr

  ******* Find switching point at most symmetric w ********
  let lowest_asym = 100
  let best_w_index = 0 ; Find most symmetric w
  let index = 0
  let tolerance = 1p ; We let the asymmetricity be plus/minus 1p of 0 

  repeat $&total_iterations 

    let asym = abs(asymmetricity[index] - 1p)
    let current_w_pmos = width[index]

    if asym < lowest_asym ; If we have something smaller, set it as the best goal and repeat
      let best_w_index = index
      let lowest_asym = asym

    end
    
    let index = index + 1
  end

  * Now that we have the best width, we now need to move towards getting the switching point

  let chosen_switching_point = switching_points[best_w_index]

end

.endc
"
