name=VARY_NMOS only_toplevel=true spice_ignore=false value="
*.options savecurrents

.control


set curplot = new
set ax = $curplot


let step_nmos=1
let step_pmos=1

let index_nmos=0
let index_pmos= 0

let final_w_nmos=11
let final_w_pmos=60

let current_w_nmos=10

let total_iterations_nmos = ceil(abs(final_w_nmos - current_w_nmos)/step_nmos)
let total_iterations_pmos = ceil(abs(final_w_pmos - current_w_pmos)/step_pmos)

let net_switching_points = vector(total_iterations_nmos)
let net_asymmetricity = vector(total_iterations_nmos)
let width_nmos = vector(total_iterations_nmos)


let switching_points = vector(total_iterations_pmos)
let asymmetricity = vector(total_iterations_pmos)
let width_pmos = vector(total_iterations_pmos)


***** Start varying nmos widths ****
while current_w_nmos < final_w_nmos
  set current_w_pmos=10

  alter m.xm1.msky130_fd_pr__nfet_01v8 W=current_w_nmos

**** Start varying pmos widths ******
  while current_w_pmos < final_w_pmos

    alter m.xm2.msky130_fd_pr__pfet_01v8 W=current_w_pmos

******* Asymmetricity simulation with pulse of 50n with 1/2 duty cycle ********
    tran 10p 50n 

    meas tran rise_time TRIG v(out) VAL=0.1 RISE=1 TARG v(out) VAL=1.62 RISE=1 
    meas tran fall_time TRIG v(out) VAL=1.62 FALL=1 TARG v(out) VAL=0.1 FALL=1

    set global_rise_fall_time = abs ( $&rise_time - $&fall_time )

    set curplot = {$ax}
    let asymmetricity[index_pmos] = $global_rise_fall_time



******* Switching point simulation ********
    dc vin 0 1.8 1m 

    meas dc switching_point WHEN v(out)=v(in) CROSS=LAST
    set global_switching_point = $&switching_point

    set curplot = {$ax}
    let switching_points[index_pmos] = $global_switching_point
    let width_pmos[index_pmos] = current_w_pmos

    let current_w_pmos = current_w_pmos + step_pmos
    let index_pmos = index_pmos + 1

  end

**** Stop varying pmos widths ******



******* Find switching point at most symmetric w (this is per nmos iteration) ********
  let lowest_asym = 100
  let best_w_index = 0 
  let iterate_pmos = 0
  let tolerance = 1p 
 * We let the asymmetricity be plus/minus 1p of 0 

  repeat $&total_iterations_pmos 

    let asym = abs({$ax}.asymmetricity[iterate_pmos] - 1p)
    let current_w_pmos = {$ax}.width_pmos[iterate_pmos]

    if asym < lowest_asym 
      let best_w_index = iterate_pmos
      let lowest_asym = asym
    end
    
    let iterate_pmos = iterate_pmos + 1
  end

* Now that we have the best width, we now need to move towards getting the switching point

* Select the cream of the crop 
  set curplot = {$ax}
  let net_switching_points[index_nmos] = {$ax}.switching_points[best_w_index]
  let net_asymmetricity[index_nmos] = {$ax}.asymmetricity[best_w_index]

* Associate it to the nmos value
  let width_nmos[index_nmos] = current_w_nmos



  let index_nmos = index_nmos + 1
  let current_w_nmos = current_w_nmos + step_nmos

end

**** Stop varying nmos widths **** 

set nolegend

******* Plot results ********
plot {$ax}.net_switching_points vs {$ax}.width_nmos
plot {$ax}.net_asymmetricity vs {$ax}.width_nmos
.endc
"
