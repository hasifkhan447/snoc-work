** sch_path: /home/hak/work/mobility.sch
**.subckt mobility
Vgs VGS GND 1.8
Vdd VDD GND 1.8
XM3 VDD net2 GND GND sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 GND net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
E1 net2 GND VOL=' V(Vgs) '
E2 VDD net1 VOL=' V(Vgs) '
**** begin user architecture code



.options savecurrents

.control
save all
*dc vgs 0 1.8 0.01 vdd 0.01 1.8 0.2
*dc vdd 0.01 1.8 0.01
dc vgs 0 1.8 0.01
let id_nmos=@m.xm3.msky130_fd_pr__nfet_01v8[id]
let id_pmos=@m.xm4.msky130_fd_pr__pfet_01v8[id]

plot deriv(sqrt(id_nmos))^2/deriv(sqrt(id_pmos))^2 title 'V_DD characteristic' xlabel 'V_DD' ylabel 'Ratio of derivatives'

write characterization.raw

set appendwrite
.endc


.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VGS
.GLOBAL VDD
.end
